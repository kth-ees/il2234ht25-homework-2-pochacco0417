module shift_register_tb;

// complete here

endmodule