module up_down_counter_tb;

// complete here

endmodule