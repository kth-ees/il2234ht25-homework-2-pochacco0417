module LFSR_6bit_tb;

// complete here

endmodule