module frequency_divider (input logic clk,
                          input logic rst_n,
                          output logic divider_out);
  
  // complete here

  endmodule