module registerfile_tb;

// complete here

endmodule