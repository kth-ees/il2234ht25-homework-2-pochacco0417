module frequency_divider_tb;

//complete here

endmodule